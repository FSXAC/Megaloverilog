// Register file is a collection of registers
// Handles incoming write and address signals

// Total of 8 registers, 3 bit address required

module RegisterFile(
	input logic [15:0] data_in,
	input logic [2:0] write_addr, read_addr,
	input 

	output logic [15:0] data_out,
)